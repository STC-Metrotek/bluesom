// soc.v

// Generated using ACDS version 14.0 200 at 2016.11.22.17:16:17

`timescale 1 ps / 1 ps
module soc (
		output wire [14:0] memory_mem_a,                     //      memory.mem_a
		output wire [2:0]  memory_mem_ba,                    //            .mem_ba
		output wire        memory_mem_ck,                    //            .mem_ck
		output wire        memory_mem_ck_n,                  //            .mem_ck_n
		output wire        memory_mem_cke,                   //            .mem_cke
		output wire        memory_mem_cs_n,                  //            .mem_cs_n
		output wire        memory_mem_ras_n,                 //            .mem_ras_n
		output wire        memory_mem_cas_n,                 //            .mem_cas_n
		output wire        memory_mem_we_n,                  //            .mem_we_n
		output wire        memory_mem_reset_n,               //            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                    //            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                   //            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                 //            .mem_dqs_n
		output wire        memory_mem_odt,                   //            .mem_odt
		output wire [3:0]  memory_mem_dm,                    //            .mem_dm
		input  wire        memory_oct_rzqin,                 //            .oct_rzqin
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,  //      hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,    //            .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,    //            .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,    //            .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,    //            .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,    //            .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,    //            .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,     //            .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,  //            .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,  //            .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,  //            .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,    //            .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,    //            .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,    //            .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,      //            .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,      //            .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,      //            .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,      //            .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,      //            .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,      //            .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,      //            .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,       //            .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,       //            .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,      //            .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,       //            .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,       //            .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,       //            .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,       //            .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,       //            .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,       //            .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,       //            .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,       //            .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,       //            .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,       //            .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,      //            .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,      //            .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,      //            .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,      //            .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,      //            .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,      //            .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,      //            .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,      //            .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO44,   //            .hps_io_gpio_inst_GPIO44
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO09, //            .hps_io_gpio_inst_LOANIO09
		input  wire        clk_25m_clk,                      //     clk_25m.clk
		output wire [66:0] hps_loan_io_in,                   // hps_loan_io.in
		input  wire [66:0] hps_loan_io_out,                  //            .out
		input  wire [66:0] hps_loan_io_oe,                   //            .oe
		input  wire        fpga_regs_waitrequest,            //   fpga_regs.waitrequest
		input  wire [31:0] fpga_regs_readdata,               //            .readdata
		input  wire        fpga_regs_readdatavalid,          //            .readdatavalid
		output wire [0:0]  fpga_regs_burstcount,             //            .burstcount
		output wire [31:0] fpga_regs_writedata,              //            .writedata
		output wire [7:0]  fpga_regs_address,                //            .address
		output wire        fpga_regs_write,                  //            .write
		output wire        fpga_regs_read,                   //            .read
		output wire [3:0]  fpga_regs_byteenable,             //            .byteenable
		output wire        fpga_regs_debugaccess,            //            .debugaccess
		output wire        clk_100m_clk                      //    clk_100m.clk
	);

	wire         hps_0_h2f_axi_master_awvalid;                          // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire   [2:0] hps_0_h2f_axi_master_arsize;                           // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire   [1:0] hps_0_h2f_axi_master_arlock;                           // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [3:0] hps_0_h2f_axi_master_awcache;                          // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire         hps_0_h2f_axi_master_arready;                          // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [11:0] hps_0_h2f_axi_master_arid;                             // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire         hps_0_h2f_axi_master_rready;                           // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire         hps_0_h2f_axi_master_bready;                           // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire   [2:0] hps_0_h2f_axi_master_awsize;                           // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire   [2:0] hps_0_h2f_axi_master_awprot;                           // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire         hps_0_h2f_axi_master_arvalid;                          // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [2:0] hps_0_h2f_axi_master_arprot;                           // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire  [11:0] hps_0_h2f_axi_master_bid;                              // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire   [3:0] hps_0_h2f_axi_master_arlen;                            // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire         hps_0_h2f_axi_master_awready;                          // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire  [11:0] hps_0_h2f_axi_master_awid;                             // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire         hps_0_h2f_axi_master_bvalid;                           // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire  [11:0] hps_0_h2f_axi_master_wid;                              // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [1:0] hps_0_h2f_axi_master_awlock;                           // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [1:0] hps_0_h2f_axi_master_awburst;                          // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [1:0] hps_0_h2f_axi_master_bresp;                            // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                            // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_rvalid;                           // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire  [31:0] hps_0_h2f_axi_master_wdata;                            // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_wready;                           // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                          // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire  [31:0] hps_0_h2f_axi_master_rdata;                            // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire  [29:0] hps_0_h2f_axi_master_araddr;                           // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [3:0] hps_0_h2f_axi_master_arcache;                          // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire   [3:0] hps_0_h2f_axi_master_awlen;                            // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                           // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire  [11:0] hps_0_h2f_axi_master_rid;                              // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_wvalid;                           // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [1:0] hps_0_h2f_axi_master_rresp;                            // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire         hps_0_h2f_axi_master_wlast;                            // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire         hps_0_h2f_axi_master_rlast;                            // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;          // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire   [9:0] mm_interconnect_0_onchip_memory_s1_address;            // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;         // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire         mm_interconnect_0_onchip_memory_s1_clken;              // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_onchip_memory_s1_write;              // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;           // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;         // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;  // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata; // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_waitrequest;          // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire   [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;           // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;            // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire   [7:0] mm_interconnect_0_mm_bridge_0_s0_address;              // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_0_mm_bridge_0_s0_write;                // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire         mm_interconnect_0_mm_bridge_0_s0_read;                 // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;             // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_debugaccess;          // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire         mm_interconnect_0_mm_bridge_0_s0_readdatavalid;        // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;           // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire  [31:0] hps_0_f2h_irq0_irq;                                    // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                    // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> pll_0:rst
	wire         hps_0_h2f_reset_reset;                                 // hps_0:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                    // rst_controller_001:reset_out -> [mm_bridge_0:reset, mm_interconnect_0:onchip_memory_reset1_reset_bridge_in_reset_reset, onchip_memory:reset, sysid_qsys_0:reset_n]

	soc_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.h2f_loan_in               (hps_loan_io_in),                   //    h2f_loan_io.in
		.h2f_loan_out              (hps_loan_io_out),                  //               .out
		.h2f_loan_oe               (hps_loan_io_oe),                   //               .oe
		.mem_a                     (memory_mem_a),                     //         memory.mem_a
		.mem_ba                    (memory_mem_ba),                    //               .mem_ba
		.mem_ck                    (memory_mem_ck),                    //               .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                  //               .mem_ck_n
		.mem_cke                   (memory_mem_cke),                   //               .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                  //               .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                 //               .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                 //               .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                  //               .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),               //               .mem_reset_n
		.mem_dq                    (memory_mem_dq),                    //               .mem_dq
		.mem_dqs                   (memory_mem_dqs),                   //               .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                 //               .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                   //               .mem_odt
		.mem_dm                    (memory_mem_dm),                    //               .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                 //               .oct_rzqin
		.hps_io_emac1_inst_TX_CLK  (hps_io_hps_io_emac1_inst_TX_CLK),  //         hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0    (hps_io_hps_io_emac1_inst_TXD0),    //               .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1    (hps_io_hps_io_emac1_inst_TXD1),    //               .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2    (hps_io_hps_io_emac1_inst_TXD2),    //               .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3    (hps_io_hps_io_emac1_inst_TXD3),    //               .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0    (hps_io_hps_io_emac1_inst_RXD0),    //               .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO    (hps_io_hps_io_emac1_inst_MDIO),    //               .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC     (hps_io_hps_io_emac1_inst_MDC),     //               .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL  (hps_io_hps_io_emac1_inst_RX_CTL),  //               .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL  (hps_io_hps_io_emac1_inst_TX_CTL),  //               .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK  (hps_io_hps_io_emac1_inst_RX_CLK),  //               .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1    (hps_io_hps_io_emac1_inst_RXD1),    //               .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2    (hps_io_hps_io_emac1_inst_RXD2),    //               .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3    (hps_io_hps_io_emac1_inst_RXD3),    //               .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0      (hps_io_hps_io_qspi_inst_IO0),      //               .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1      (hps_io_hps_io_qspi_inst_IO1),      //               .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2      (hps_io_hps_io_qspi_inst_IO2),      //               .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3      (hps_io_hps_io_qspi_inst_IO3),      //               .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0      (hps_io_hps_io_qspi_inst_SS0),      //               .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK      (hps_io_hps_io_qspi_inst_CLK),      //               .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD      (hps_io_hps_io_sdio_inst_CMD),      //               .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0       (hps_io_hps_io_sdio_inst_D0),       //               .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1       (hps_io_hps_io_sdio_inst_D1),       //               .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK      (hps_io_hps_io_sdio_inst_CLK),      //               .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2       (hps_io_hps_io_sdio_inst_D2),       //               .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3       (hps_io_hps_io_sdio_inst_D3),       //               .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0       (hps_io_hps_io_usb1_inst_D0),       //               .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1       (hps_io_hps_io_usb1_inst_D1),       //               .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2       (hps_io_hps_io_usb1_inst_D2),       //               .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3       (hps_io_hps_io_usb1_inst_D3),       //               .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4       (hps_io_hps_io_usb1_inst_D4),       //               .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5       (hps_io_hps_io_usb1_inst_D5),       //               .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6       (hps_io_hps_io_usb1_inst_D6),       //               .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7       (hps_io_hps_io_usb1_inst_D7),       //               .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK      (hps_io_hps_io_usb1_inst_CLK),      //               .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP      (hps_io_hps_io_usb1_inst_STP),      //               .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR      (hps_io_hps_io_usb1_inst_DIR),      //               .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT      (hps_io_hps_io_usb1_inst_NXT),      //               .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX      (hps_io_hps_io_uart0_inst_RX),      //               .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX      (hps_io_hps_io_uart0_inst_TX),      //               .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA      (hps_io_hps_io_i2c0_inst_SDA),      //               .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL      (hps_io_hps_io_i2c0_inst_SCL),      //               .hps_io_i2c0_inst_SCL
		.hps_io_gpio_inst_GPIO44   (hps_io_hps_io_gpio_inst_GPIO44),   //               .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_LOANIO09 (hps_io_hps_io_gpio_inst_LOANIO09), //               .hps_io_gpio_inst_LOANIO09
		.h2f_rst_n                 (hps_0_h2f_reset_reset),            //      h2f_reset.reset_n
		.h2f_axi_clk               (clk_100m_clk),                     //  h2f_axi_clock.clk
		.h2f_AWID                  (hps_0_h2f_axi_master_awid),        // h2f_axi_master.awid
		.h2f_AWADDR                (hps_0_h2f_axi_master_awaddr),      //               .awaddr
		.h2f_AWLEN                 (hps_0_h2f_axi_master_awlen),       //               .awlen
		.h2f_AWSIZE                (hps_0_h2f_axi_master_awsize),      //               .awsize
		.h2f_AWBURST               (hps_0_h2f_axi_master_awburst),     //               .awburst
		.h2f_AWLOCK                (hps_0_h2f_axi_master_awlock),      //               .awlock
		.h2f_AWCACHE               (hps_0_h2f_axi_master_awcache),     //               .awcache
		.h2f_AWPROT                (hps_0_h2f_axi_master_awprot),      //               .awprot
		.h2f_AWVALID               (hps_0_h2f_axi_master_awvalid),     //               .awvalid
		.h2f_AWREADY               (hps_0_h2f_axi_master_awready),     //               .awready
		.h2f_WID                   (hps_0_h2f_axi_master_wid),         //               .wid
		.h2f_WDATA                 (hps_0_h2f_axi_master_wdata),       //               .wdata
		.h2f_WSTRB                 (hps_0_h2f_axi_master_wstrb),       //               .wstrb
		.h2f_WLAST                 (hps_0_h2f_axi_master_wlast),       //               .wlast
		.h2f_WVALID                (hps_0_h2f_axi_master_wvalid),      //               .wvalid
		.h2f_WREADY                (hps_0_h2f_axi_master_wready),      //               .wready
		.h2f_BID                   (hps_0_h2f_axi_master_bid),         //               .bid
		.h2f_BRESP                 (hps_0_h2f_axi_master_bresp),       //               .bresp
		.h2f_BVALID                (hps_0_h2f_axi_master_bvalid),      //               .bvalid
		.h2f_BREADY                (hps_0_h2f_axi_master_bready),      //               .bready
		.h2f_ARID                  (hps_0_h2f_axi_master_arid),        //               .arid
		.h2f_ARADDR                (hps_0_h2f_axi_master_araddr),      //               .araddr
		.h2f_ARLEN                 (hps_0_h2f_axi_master_arlen),       //               .arlen
		.h2f_ARSIZE                (hps_0_h2f_axi_master_arsize),      //               .arsize
		.h2f_ARBURST               (hps_0_h2f_axi_master_arburst),     //               .arburst
		.h2f_ARLOCK                (hps_0_h2f_axi_master_arlock),      //               .arlock
		.h2f_ARCACHE               (hps_0_h2f_axi_master_arcache),     //               .arcache
		.h2f_ARPROT                (hps_0_h2f_axi_master_arprot),      //               .arprot
		.h2f_ARVALID               (hps_0_h2f_axi_master_arvalid),     //               .arvalid
		.h2f_ARREADY               (hps_0_h2f_axi_master_arready),     //               .arready
		.h2f_RID                   (hps_0_h2f_axi_master_rid),         //               .rid
		.h2f_RDATA                 (hps_0_h2f_axi_master_rdata),       //               .rdata
		.h2f_RRESP                 (hps_0_h2f_axi_master_rresp),       //               .rresp
		.h2f_RLAST                 (hps_0_h2f_axi_master_rlast),       //               .rlast
		.h2f_RVALID                (hps_0_h2f_axi_master_rvalid),      //               .rvalid
		.h2f_RREADY                (hps_0_h2f_axi_master_rready),      //               .rready
		.f2h_irq_p0                (hps_0_f2h_irq0_irq),               //       f2h_irq0.irq
		.f2h_irq_p1                (hps_0_f2h_irq1_irq)                //       f2h_irq1.irq
	);

	soc_pll_0 pll_0 (
		.refclk   (clk_25m_clk),                    //  refclk.clk
		.rst      (rst_controller_reset_out_reset), //   reset.reset
		.outclk_0 (clk_100m_clk),                   // outclk0.clk
		.locked   ()                                // (terminated)
	);

	soc_onchip_memory onchip_memory (
		.clk        (clk_100m_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (1'b0)                                           // (terminated)
	);

	soc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_100m_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (8),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_100m_clk),                                   //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (fpga_regs_waitrequest),                          //    m0.waitrequest
		.m0_readdata      (fpga_regs_readdata),                             //      .readdata
		.m0_readdatavalid (fpga_regs_readdatavalid),                        //      .readdatavalid
		.m0_burstcount    (fpga_regs_burstcount),                           //      .burstcount
		.m0_writedata     (fpga_regs_writedata),                            //      .writedata
		.m0_address       (fpga_regs_address),                              //      .address
		.m0_write         (fpga_regs_write),                                //      .write
		.m0_read          (fpga_regs_read),                                 //      .read
		.m0_byteenable    (fpga_regs_byteenable),                           //      .byteenable
		.m0_debugaccess   (fpga_regs_debugaccess)                           //      .debugaccess
	);

	soc_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                        (hps_0_h2f_axi_master_awid),                             //                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                      (hps_0_h2f_axi_master_awaddr),                           //                                           .awaddr
		.hps_0_h2f_axi_master_awlen                       (hps_0_h2f_axi_master_awlen),                            //                                           .awlen
		.hps_0_h2f_axi_master_awsize                      (hps_0_h2f_axi_master_awsize),                           //                                           .awsize
		.hps_0_h2f_axi_master_awburst                     (hps_0_h2f_axi_master_awburst),                          //                                           .awburst
		.hps_0_h2f_axi_master_awlock                      (hps_0_h2f_axi_master_awlock),                           //                                           .awlock
		.hps_0_h2f_axi_master_awcache                     (hps_0_h2f_axi_master_awcache),                          //                                           .awcache
		.hps_0_h2f_axi_master_awprot                      (hps_0_h2f_axi_master_awprot),                           //                                           .awprot
		.hps_0_h2f_axi_master_awvalid                     (hps_0_h2f_axi_master_awvalid),                          //                                           .awvalid
		.hps_0_h2f_axi_master_awready                     (hps_0_h2f_axi_master_awready),                          //                                           .awready
		.hps_0_h2f_axi_master_wid                         (hps_0_h2f_axi_master_wid),                              //                                           .wid
		.hps_0_h2f_axi_master_wdata                       (hps_0_h2f_axi_master_wdata),                            //                                           .wdata
		.hps_0_h2f_axi_master_wstrb                       (hps_0_h2f_axi_master_wstrb),                            //                                           .wstrb
		.hps_0_h2f_axi_master_wlast                       (hps_0_h2f_axi_master_wlast),                            //                                           .wlast
		.hps_0_h2f_axi_master_wvalid                      (hps_0_h2f_axi_master_wvalid),                           //                                           .wvalid
		.hps_0_h2f_axi_master_wready                      (hps_0_h2f_axi_master_wready),                           //                                           .wready
		.hps_0_h2f_axi_master_bid                         (hps_0_h2f_axi_master_bid),                              //                                           .bid
		.hps_0_h2f_axi_master_bresp                       (hps_0_h2f_axi_master_bresp),                            //                                           .bresp
		.hps_0_h2f_axi_master_bvalid                      (hps_0_h2f_axi_master_bvalid),                           //                                           .bvalid
		.hps_0_h2f_axi_master_bready                      (hps_0_h2f_axi_master_bready),                           //                                           .bready
		.hps_0_h2f_axi_master_arid                        (hps_0_h2f_axi_master_arid),                             //                                           .arid
		.hps_0_h2f_axi_master_araddr                      (hps_0_h2f_axi_master_araddr),                           //                                           .araddr
		.hps_0_h2f_axi_master_arlen                       (hps_0_h2f_axi_master_arlen),                            //                                           .arlen
		.hps_0_h2f_axi_master_arsize                      (hps_0_h2f_axi_master_arsize),                           //                                           .arsize
		.hps_0_h2f_axi_master_arburst                     (hps_0_h2f_axi_master_arburst),                          //                                           .arburst
		.hps_0_h2f_axi_master_arlock                      (hps_0_h2f_axi_master_arlock),                           //                                           .arlock
		.hps_0_h2f_axi_master_arcache                     (hps_0_h2f_axi_master_arcache),                          //                                           .arcache
		.hps_0_h2f_axi_master_arprot                      (hps_0_h2f_axi_master_arprot),                           //                                           .arprot
		.hps_0_h2f_axi_master_arvalid                     (hps_0_h2f_axi_master_arvalid),                          //                                           .arvalid
		.hps_0_h2f_axi_master_arready                     (hps_0_h2f_axi_master_arready),                          //                                           .arready
		.hps_0_h2f_axi_master_rid                         (hps_0_h2f_axi_master_rid),                              //                                           .rid
		.hps_0_h2f_axi_master_rdata                       (hps_0_h2f_axi_master_rdata),                            //                                           .rdata
		.hps_0_h2f_axi_master_rresp                       (hps_0_h2f_axi_master_rresp),                            //                                           .rresp
		.hps_0_h2f_axi_master_rlast                       (hps_0_h2f_axi_master_rlast),                            //                                           .rlast
		.hps_0_h2f_axi_master_rvalid                      (hps_0_h2f_axi_master_rvalid),                           //                                           .rvalid
		.hps_0_h2f_axi_master_rready                      (hps_0_h2f_axi_master_rready),                           //                                           .rready
		.pll_0_outclk0_clk                                (clk_100m_clk),                                          //                              pll_0_outclk0.clk
		.onchip_memory_reset1_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // onchip_memory_reset1_reset_bridge_in_reset.reset
		.mm_bridge_0_s0_address                           (mm_interconnect_0_mm_bridge_0_s0_address),              //                             mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                             (mm_interconnect_0_mm_bridge_0_s0_write),                //                                           .write
		.mm_bridge_0_s0_read                              (mm_interconnect_0_mm_bridge_0_s0_read),                 //                                           .read
		.mm_bridge_0_s0_readdata                          (mm_interconnect_0_mm_bridge_0_s0_readdata),             //                                           .readdata
		.mm_bridge_0_s0_writedata                         (mm_interconnect_0_mm_bridge_0_s0_writedata),            //                                           .writedata
		.mm_bridge_0_s0_burstcount                        (mm_interconnect_0_mm_bridge_0_s0_burstcount),           //                                           .burstcount
		.mm_bridge_0_s0_byteenable                        (mm_interconnect_0_mm_bridge_0_s0_byteenable),           //                                           .byteenable
		.mm_bridge_0_s0_readdatavalid                     (mm_interconnect_0_mm_bridge_0_s0_readdatavalid),        //                                           .readdatavalid
		.mm_bridge_0_s0_waitrequest                       (mm_interconnect_0_mm_bridge_0_s0_waitrequest),          //                                           .waitrequest
		.mm_bridge_0_s0_debugaccess                       (mm_interconnect_0_mm_bridge_0_s0_debugaccess),          //                                           .debugaccess
		.onchip_memory_s1_address                         (mm_interconnect_0_onchip_memory_s1_address),            //                           onchip_memory_s1.address
		.onchip_memory_s1_write                           (mm_interconnect_0_onchip_memory_s1_write),              //                                           .write
		.onchip_memory_s1_readdata                        (mm_interconnect_0_onchip_memory_s1_readdata),           //                                           .readdata
		.onchip_memory_s1_writedata                       (mm_interconnect_0_onchip_memory_s1_writedata),          //                                           .writedata
		.onchip_memory_s1_byteenable                      (mm_interconnect_0_onchip_memory_s1_byteenable),         //                                           .byteenable
		.onchip_memory_s1_chipselect                      (mm_interconnect_0_onchip_memory_s1_chipselect),         //                                           .chipselect
		.onchip_memory_s1_clken                           (mm_interconnect_0_onchip_memory_s1_clken),              //                                           .clken
		.sysid_qsys_0_control_slave_address               (mm_interconnect_0_sysid_qsys_0_control_slave_address),  //                 sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata              (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)  //                                           .readdata
	);

	soc_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (clk_25m_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_100m_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
